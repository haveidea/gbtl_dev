// single_adder.v

// Generated using ACDS version 16.1 196

`timescale 1 ps / 1 ps
module single_adder (
                input  wire [1:0]  aclr,   //   aclr.aclr
                input  wire [31:0] ax,     //     ax.ax
                input  wire [31:0] ay,     //     ay.ay
                output wire [31:0] result  // result.result
        );
//`ifndef SIMU
        single_adder_comb   fpdsp_block_0 (
                .aclr   (aclr),   //   aclr.aclr
                .result (result), // result.result
                .ax     (ax),     //     ax.ax
                .ay     (ay)      //     ay.ay
        );
//`else
// DW_fp_add fp_adder(.a(ax), .b(ay), .rnd(3'b000), .z(result), .status());
//`endif

endmodule
