//
//---------------------------------------------------------------------------
// LiM memory block for segment for both buffer and stage output
//  
//  
//---------------------------------------------------------------------------
//
`include "definitions.vh"

module segment_memory_reg #(
   parameter
     NUM_BUFF_SO_WORDS_SEG = `NUM_BUFF_SO_WORDS_SEG,	   
     DATA_WIDTH = `DATA_WIDTH_BUFF_SO_SEG,
     BITS_ADDR_SEG = `BITS_ADDR_SEG) (

   input rst_b, clk, wr_en, mandatory_bubble,
   input [BITS_ADDR_SEG - 1 : 0] rd_addr_seg, 
   input [BITS_ADDR_SEG - 1 : 0] adv_wr_addr_seg,  
   input [DATA_WIDTH - 1 : 0] data_in_buff, data_in_so,
							  
   output logic [DATA_WIDTH - 1 : 0] dout_buff, dout_so);

//reg memory
//valiables with unpacked are not displayed in NCSim simulation, but works fine   
logic [NUM_BUFF_SO_WORDS_SEG - 1 : 0] [DATA_WIDTH - 1 : 0] buff_reg;   
logic [NUM_BUFF_SO_WORDS_SEG - 1 : 0] [DATA_WIDTH - 1 : 0] so_reg;

integer i; 
always_ff @(posedge clk) begin    
   if(~rst_b) begin
      for (i = 0; i < NUM_BUFF_SO_WORDS_SEG; i = i + 1) begin
	 buff_reg[i] <=  0; 
	 so_reg[i] <=  0;
      end
   end
   //write
   else if(wr_en && rst_b) begin
      buff_reg[adv_wr_addr_seg] <= data_in_buff;
      so_reg[adv_wr_addr_seg] <= data_in_so;
   end
end   

//this is for nonpipelined version. technically this will functionally work for pipelined version too   
//assign dout_buff = buff_reg[rd_addr_seg];
//assign dout_so = so_reg[rd_addr_seg];

//this is for pipelined version
register #(.WIDTH(DATA_WIDTH)) reg_dout_buff(.q(dout_buff), .d(buff_reg[rd_addr_seg]), .clk, .enable(mandatory_bubble), .rst_b(rst_b));
register #(.WIDTH(DATA_WIDTH)) reg_dout_so(.q(dout_so), .d(so_reg[rd_addr_seg]), .clk, .enable(mandatory_bubble), .rst_b(rst_b));   
   

//********** INPUT FLOPS **********  
/*
integer i;
always_ff @ (posedge clk) begin
   if(~rst_b) begin
      for (i = 0; i < NUM_BUFF_SO_WORDS_SEG; i = i + 1) begin
	 buff_reg[i] <=  0; 
	 so_reg[i] <=  0;
      end
   end
   else begin
      for (i = 0; i < NUM_BUFF_SO_WORDS_SEG; i = i + 1) begin
	 buff_reg[i] <= decoded_reg_type_mem[i] ? data_in_buff : buff_reg[i]; //even though writing, we use rd wl in WORK mode
	 so_reg[i] <= decoded_reg_type_mem[i] ? data_in_so : so_reg[i];// as we need wl ready before clk edge. This is because FLOP is generated by the tool. After the clock edge, whatever wordline is active immediately, data will be written to that. We activate the wordlines in the same cycle where data is written. For registers, it will not allow the time needed to activate the wordlines from address. So the data may get corrupted for registers. For LiM, this is not an issue as it acts as a black box and wordline activation delay and data write is taken care of internally. For read, this issue is not a problem for registers either. Because for registers, read process doesn't have to be flopped and corruption cannot happen. In the worst case, data will show up at the BLs late because of the wordline activation delay. 
      end
   end
end
*/
endmodule

